--- top level entity
library ieee;
use ieee.std_logic_1164.all;
use iee.numeric_std.all

library work;
use control_generic_pkg.all